module demux_tb ();
	