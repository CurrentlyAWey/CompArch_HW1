module delay(
	input d,
	output q);